module riscv_soft_d_cache(
			  clk,
			  reset,
			  req_ready,
			  req_valid,
			  req_op,
			  req_op_type,
			  req_addr,
			  req_data,
			  resp_valid,
			  resp_data
			  );


endmodule // riscv_soft_d_cache
