module riscv_soft_i_cache(
			  clk,
			  reset,
			  req_ready,
			  req_valid,
			  req_addr,
			  resp_valid,
			  resp_data
			  );


endmodule // riscv_soft_i_cache
